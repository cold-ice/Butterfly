LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY mult_add_tb IS

--PORT();

END mult_add_tb;


ARCHITECTURE behavioural OF mult_add_tb IS

COMPONENT ADDER
PORT(	DATA_IN0	: IN SIGNED(30 downto 0):=(others=>'0');
	DATA_IN1	: IN SIGNED(30 downto 0):=(others=>'0');
	C0		: IN STD_LOGIC:='0';
	DATA_OUT	: OUT SIGNED(30 downto 0):=(others=>'0')
);
END COMPONENT;

COMPONENT MULTIPLIER
PORT(	DATA_IN0	: IN SIGNED(15 downto 0):=(others=>'0');
	DATA_IN1	: IN SIGNED(15 downto 0):=(others=>'0');
	DATA_OUT	: OUT SIGNED(31 downto 0):=(others=>'0')
);
END COMPONENT;

COMPONENT SHIFTER_X2
PORT(	DATA_IN		: IN SIGNED(15 downto 0):=(others=>'0');
	DATA_OUT	: OUT SIGNED(15 downto 0):=(others=>'0')
);
END COMPONENT;

SIGNAL DATA_IN0, DATA_IN1 : SIGNED(30 downto 0);
SIGNAL C0 : STD_LOGIC;

BEGIN

add: ADDER		PORT MAP(DATA_IN0, DATA_IN1, C0);
mult: MULTIPLIER	PORT MAP(DATA_IN0(30 downto 15), DATA_IN1(30 downto 15));
shf: SHIFTER_X2		PORT MAP(DATA_IN0(30 downto 15));

signals: PROCESS
BEGIN
DATA_IN0<="0000000000000001000000000000000";
DATA_IN1<="0000000000000001100000000000000";
C0<='0';
wait for 40 ns;
DATA_IN0<="1111111111111110111111111111111"; -- -32769
DATA_IN1<="1111111111111110000000000000000"; -- -65536
C0<='0';
wait for 40 ns;
DATA_IN0<="0000000000000001000000000000000";
DATA_IN1<="1111111111111111000000000000000";
C0<='0';
wait for 40 ns;
DATA_IN0<="0000000000000001000000000000000";
DATA_IN1<="0000000000000001100000000000000";
C0<='1';
wait for 40 ns;
DATA_IN0<="1111111111111110111111111111111";
DATA_IN1<="1111111111111110000000000000000";
C0<='1';
wait for 40 ns;
DATA_IN0<="0000000000000001000000000000000";
DATA_IN1<="1111111111111111000000000000000";
C0<='1';
wait for 40 ns;
END PROCESS;

END behavioural;