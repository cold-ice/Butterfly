library IEEE;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY REG2 IS
GENERIC (SIZE			: INTEGER);
PORT(		CLOCK		 	: IN STD_LOGIC;
			ENABLE		: IN STD_LOGIC;
			CLEAR			: IN STD_LOGIC;
			INPUT			: IN STD_LOGIC_VECTOR(SIZE downto 0);
			OUTPUT		: OUT STD_LOGIC_VECTOR(SIZE downto 0)
);
END ENTITY;

ARCHITECTURE behavioural OF REG2 IS

BEGIN

FF: PROCESS(CLOCK, CLEAR)
BEGIN
IF(CLEAR = '1') THEN
	OUTPUT<= (others =>'0');
ELSIF(RISING_EDGE(CLOCK)) THEN
	IF(ENABLE = '1') THEN
		OUTPUT <= INPUT;
	END IF;
END IF;
END PROCESS;

END behavioural;