LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY ROUNDER_tb IS

--PORT();

END ROUNDER_tb;


ARCHITECTURE behavioural OF ROUNDER_tb IS

COMPONENT ROUNDER
PORT(	DATA_IN	: IN SIGNED(30 downto 0):=(others=>'0');
		DATA_OUT	: OUT SIGNED(15 downto 0):=(others=>'0')
);
END COMPONENT;

SIGNAL DATA_IN : SIGNED(30 downto 0);

BEGIN

ROUND: ROUNDER	PORT MAP(DATA_IN);

signals: PROCESS
BEGIN
DATA_IN<="0000000000000000"&"100000000000000"; --NO
wait for 40 ns;
DATA_IN<="0000000000000000"&"100000000000001"; --YES
wait for 40 ns;
DATA_IN<="0000000000000001"&"100000000000000"; --YES
wait for 40 ns;
DATA_IN<="1000000000000010"&"100000000000000"; --NO
wait for 40 ns;
DATA_IN<="1000000000000010"&"100000000000001"; --YES
wait for 40 ns;
DATA_IN<="1000000000000011"&"100000000000000"; --YES
wait for 40 ns;
wait;
END PROCESS;

END behavioural;